module add4bit_hdl (
    input   logic   
);

endmodule