module seg7animation