module test_mux7seg (
    input   logic       clk,
    input
);
    
endmodule