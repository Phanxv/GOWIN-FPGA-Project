module simple_io(
    input logic tws0,
    output logic led0
);

    assign led0 = tws0;

endmodule : simple_io